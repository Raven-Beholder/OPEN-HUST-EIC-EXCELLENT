module  decoder3_8(//3_8????
      input [2:0] A,//????a,[2:0]????
      input g1,
      input g2,
      input g3,//????1~3
      output reg[7:0] y//????y?[7:0]????
      );

always @(*) begin
        if({g1,g2,g3} != 3'b100) //g1 g2 g3??????????100???(????)
           y <= 8'h00;
        else 
           case(A)
              3'b000: y <= 8'b0000_0001; 
              3'b001: y <= 8'b0000_0010; 
              3'b010: y <= 8'b0000_0100; 
              3'b011: y <= 8'b0000_1000; 
              3'b100: y <= 8'b0001_0000; 
              3'b101: y <= 8'b0010_0000; 
              3'b110: y <= 8'b0100_0000; 
              3'b111: y <= 8'b1000_0000; 
           endcase
end
endmodule