`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/03/10 15:27:19
// Design Name: 
// Module Name:                                                              
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module decoder_4_16(
    input clk,
    input [3:0] Y,
    input rst_n,
    output reg [15:0] Q
    );
    
    
    always @(posedge clk)
        if (rst_n)
            Q <= 16'h0000;
        else
            case ({Y[3],Y[2],Y[1],Y[0]})
            4'b0000  : Q <= 16'b0000000000000001;
            4'b0001  : Q <= 16'b0000000000000010;
            4'b0010  : Q <= 16'b0000000000000100;
            4'b0011  : Q <= 16'b0000000000001000;
            4'b0100  : Q <= 16'b0000000000010000;
            4'b0101  : Q <= 16'b0000000000100000;
            4'b0110  : Q <= 16'b0000000001000000;
            4'b0111  : Q <= 16'b0000000010000000;
            4'b1000  : Q <= 16'b0000000100000000;
            4'b1001  : Q <= 16'b0000001000000000;
            4'b1010  : Q <= 16'b0000010000000000;
            4'b1011  : Q <= 16'b0000100000000000;
            4'b1100  : Q <= 16'b0001000000000000;
            4'b1101  : Q <= 16'b0010000000000000;
            4'b1110  : Q <= 16'b0100000000000000;
            4'b1111  : Q <= 16'b1000000000000000;
            default : Q <= 16'b0000000000000000;
        endcase
endmodule
